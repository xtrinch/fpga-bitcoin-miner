`timescale 1ns/1ps

// A quick define to help index 32-bit words inside a larger register.
`define IDX(x) (((x)+1)*(32)-1):((x)*(32))

// Perform a SHA-256 transformation on the given 512-bit data, and 256-bit
// initial state,
// Outputs one 256-bit hash every LOOP cycle(s).
//
// The LOOP parameter determines both the size and speed of this module.
// A value of 1 implies a fully unrolled SHA-256 calculation spanning 64 round
// modules and calculating a full SHA-256 hash every clock cycle. A value of
// 2 implies a half-unrolled loop, with 32 round modules and calculating
// a full hash in 2 clock cycles. And so forth.
module sha256_transform #(
	parameter LOOP = 6'd4
) (
	input clk,
	input feedback, // On the first count (cnt==0), load data from previous stage (feedback=0),
					// on 1..LOOP-1, take feedback from current stage (feedback=1)
	input [5:0] cnt, // where in the LOOP are we
	input [255:0] rx_state, // initial compression state
	input [511:0] rx_input, // data we'd like to hash
	output reg [255:0] tx_hash // 255 bit hash output
);
	// 64 Constants defined by the SHA-2 standard. - sqrt3(primes)
	localparam Ks = {
		32'h428a2f98, 32'h71374491, 32'hb5c0fbcf, 32'he9b5dba5,
		32'h3956c25b, 32'h59f111f1, 32'h923f82a4, 32'hab1c5ed5,
		32'hd807aa98, 32'h12835b01, 32'h243185be, 32'h550c7dc3,
		32'h72be5d74, 32'h80deb1fe, 32'h9bdc06a7, 32'hc19bf174,
		32'he49b69c1, 32'hefbe4786, 32'h0fc19dc6, 32'h240ca1cc,
		32'h2de92c6f, 32'h4a7484aa, 32'h5cb0a9dc, 32'h76f988da,
		32'h983e5152, 32'ha831c66d, 32'hb00327c8, 32'hbf597fc7,
		32'hc6e00bf3, 32'hd5a79147, 32'h06ca6351, 32'h14292967,
		32'h27b70a85, 32'h2e1b2138, 32'h4d2c6dfc, 32'h53380d13,
		32'h650a7354, 32'h766a0abb, 32'h81c2c92e, 32'h92722c85,
		32'ha2bfe8a1, 32'ha81a664b, 32'hc24b8b70, 32'hc76c51a3,
		32'hd192e819, 32'hd6990624, 32'hf40e3585, 32'h106aa070,
		32'h19a4c116, 32'h1e376c08, 32'h2748774c, 32'h34b0bcb5,
		32'h391c0cb3, 32'h4ed8aa4a, 32'h5b9cca4f, 32'h682e6ff3,
		32'h748f82ee, 32'h78a5636f, 32'h84c87814, 32'h8cc70208,
		32'h90befffa, 32'ha4506ceb, 32'hbef9a3f7, 32'hc67178f2};

	// generate the message schedule pipeline - 64 words (word is 32 bytes)
	genvar i;
	generate
		for (i = 0; i < 64/LOOP; i = i + 1) begin: HASHERS
			wire [511:0] W; // message schedule word
			wire [255:0] state; // compression state

			if(i == 0)
				sha256_digester U (
					.clk(clk), // clock
					.k(Ks[32*(63-cnt) +: 32]), // constant
					.rx_w(feedback ? W : rx_input), // if feedback use the current message schedule word, otherwise take a new one
					.rx_state(feedback ? state : rx_state), // input state, if feedback we use the state we just calculated and do not advance the pipeline
					.tx_w(W),
					.tx_state(state) // output state
				);
			else
				sha256_digester U (
					.clk(clk), // clock
					.k(Ks[32*(63-LOOP*i-cnt) +: 32]), // constant
					.rx_w(feedback ? W : HASHERS[i-1].W),
					.rx_state(feedback ? state : HASHERS[i-1].state), // input state
					.tx_w(W),
					.tx_state(state) // output state
				);
		end
	endgenerate

	// output the computed hash, it will be in the last state of the pipeline, 
	// add in the initial receiving state as per sha256
	always @ (posedge clk)
	begin
		if (!feedback) // cnt == 0
		begin
			tx_hash[`IDX(0)] <= rx_state[`IDX(0)] + HASHERS[64/LOOP-6'd1].state[`IDX(0)];
			tx_hash[`IDX(1)] <= rx_state[`IDX(1)] + HASHERS[64/LOOP-6'd1].state[`IDX(1)];
			tx_hash[`IDX(2)] <= rx_state[`IDX(2)] + HASHERS[64/LOOP-6'd1].state[`IDX(2)];
			tx_hash[`IDX(3)] <= rx_state[`IDX(3)] + HASHERS[64/LOOP-6'd1].state[`IDX(3)];
			tx_hash[`IDX(4)] <= rx_state[`IDX(4)] + HASHERS[64/LOOP-6'd1].state[`IDX(4)];
			tx_hash[`IDX(5)] <= rx_state[`IDX(5)] + HASHERS[64/LOOP-6'd1].state[`IDX(5)];
			tx_hash[`IDX(6)] <= rx_state[`IDX(6)] + HASHERS[64/LOOP-6'd1].state[`IDX(6)];
			tx_hash[`IDX(7)] <= rx_state[`IDX(7)] + HASHERS[64/LOOP-6'd1].state[`IDX(7)];
		end
	end
endmodule

module sha256_digester (
	input clk, // clock
	input [31:0] k, // constant
	input [511:0] rx_w, // message schedule, 16 words
	input [255:0] rx_state, // input state of stage (prev state)
	output reg [511:0] tx_w, // next stage of the message schedule
	output reg [255:0] tx_state // calculated next state of compression stage
);
	// temporary words declaration for use in below calculations
	wire [31:0] e0_w, e1_w, ch_w, maj_w, s0_w, s1_w;

	// new message schedule word calculation
	s0	s0_blk	(rx_w[63:32], s0_w);
	s1	s1_blk	(rx_w[479:448], s1_w);
	
	// new message schedule word
	wire [31:0] new_w = s1_w + rx_w[319:288] + s0_w + rx_w[31:0];

	// T1 and T2 reg calculation
	e0	e0_blk	(rx_state[`IDX(0)], e0_w);
	e1	e1_blk	(rx_state[`IDX(4)], e1_w);
	ch	ch_blk	(rx_state[`IDX(4)], rx_state[`IDX(5)], rx_state[`IDX(6)], ch_w);
	maj	maj_blk	(rx_state[`IDX(0)], rx_state[`IDX(1)], rx_state[`IDX(2)], maj_w);

	wire [31:0] t1 = rx_state[`IDX(7)] + e1_w + ch_w + rx_w[31:0] + k; // T1 for the compression
	wire [31:0] t2 = e0_w + maj_w; // T2 for the compression

	always @ (posedge clk)
	begin
		tx_w[511:480] <= new_w; // slide in from the left the new word of the message schedule 
		tx_w[479:0] <= rx_w[511:32]; // right shift by 1 word (32 bits)

		tx_state[`IDX(7)] <= rx_state[`IDX(6)]; // shift them all up by one word
		tx_state[`IDX(6)] <= rx_state[`IDX(5)];
		tx_state[`IDX(5)] <= rx_state[`IDX(4)];
		tx_state[`IDX(4)] <= rx_state[`IDX(3)] + t1;
		tx_state[`IDX(3)] <= rx_state[`IDX(2)];
		tx_state[`IDX(2)] <= rx_state[`IDX(1)];
		tx_state[`IDX(1)] <= rx_state[`IDX(0)];
		tx_state[`IDX(0)] <= t1 + t2;
	end
endmodule